module DE10Lite_MLP (

	///////// Clocks /////////
	input             MAX10_CLK1_50,
	
	///////// KEY /////////
	input    [1: 0]   KEY,
	
	///////// SW /////////
	input    [9: 0]   SW,
	
	///////// LEDR /////////
	output   [ 9: 0]  LEDR,
	
	///////// HEX /////////
	output   [7: 0]   HEX0,
	output   [7: 0]   HEX1,
	output   [7: 0]   HEX2,
	output   [7: 0]   HEX3,
	output   [7: 0]   HEX4,
	output   [7: 0]   HEX5,
	
	///////// SDRAM /////////
	output            DRAM_CLK,
	output            DRAM_CKE,
	output   [12: 0]  DRAM_ADDR,
	output   [ 1: 0]  DRAM_BA,
	inout    [15: 0]  DRAM_DQ,
	output            DRAM_LDQM,
	output            DRAM_UDQM,
	output            DRAM_CS_N,
	output            DRAM_WE_N,
	output            DRAM_CAS_N,
	output            DRAM_RAS_N
	);



//=======================================================
//  REG/WIRE declarations
//=======================================================

wire			[31: 0]	hex3_hex0;
wire			[15: 0]	hex5_hex4;

assign HEX0 = ~hex3_hex0[ 7: 0];
assign HEX1 = ~hex3_hex0[15: 8];
assign HEX2 = ~hex3_hex0[23:16];
assign HEX3 = ~hex3_hex0[31:24];
assign HEX4 = ~hex5_hex4[ 7: 0];
assign HEX5 = ~hex5_hex4[15: 8];


//=======================================================
//  Structural coding
//=======================================================

DE10Lite_MLP_Computer_QSYS computer_inst0 (
	
	   .clk_clk                           		(MAX10_CLK1_50),                           
		.reset_reset_n                     		(1'b1),                     
	 
		.key_external_connection_export   		(KEY),    
		.sliders_external_connection_export   	(SW),   
      .hex3_hex0_external_connection_export 	(hex3_hex0), 
      .hex5_hex4_external_connection_export 	(hex5_hex4),
		.ledr_external_connection_export 		(LEDR),
	
		//SDRAM
		.clk_sdram_clk									(DRAM_CLK),                  
		.sdram_wire_addr								(DRAM_ADDR),                
		.sdram_wire_ba									(DRAM_BA),                  
		.sdram_wire_cas_n								(DRAM_CAS_N),               
		.sdram_wire_cke								(DRAM_CKE),                 
		.sdram_wire_cs_n								(DRAM_CS_N),                
		.sdram_wire_dq									(DRAM_DQ),                  
		.sdram_wire_dqm								({DRAM_UDQM,DRAM_LDQM}),               
		.sdram_wire_ras_n								(DRAM_RAS_N),               
		.sdram_wire_we_n								(DRAM_WE_N)                 

);


endmodule
